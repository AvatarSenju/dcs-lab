----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 10/20/2018 02:57:38 PM
-- Design Name: 
-- Module Name: dff_R - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity dff_R is
    Port ( d : in STD_LOGIC;
           clk : in STD_LOGIC;
           res : in STD_LOGIC;
           q : out STD_LOGIC);
end dff_R;

architecture Behavioral of dff_R is

begin

process(d,clk,res)
begin
   if(res='1')then
        q<='0';
   else
         if(falling_edge(clk))then
             q<=d;
         end if;
   end if;
end process;

end Behavioral;
